library IEEE;
USE ieee.std_logic_1164.all;

ENTITY TripleDES IS
PORT(
	encrypt: in std_logic;
	ready: out std_logic
);
END TripleDES;

architecture comportamento of TripleDES is  
begin
end comportamento;