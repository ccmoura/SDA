ENTITY manchester is
PORT (
	A, B, Cin : in bit;
	S, Cout : out bit
);
END manchester;
architecture comportamento of manchester is 
BEGIN 
	S <= A xor B xor Cin;
	Cout <= (A and b) or (Cin and (A xor B));
END comportamento;

--somador manchester ^
--somador 32 bits v
ENTITY Somador32Bits is 
PORT (
	A : in bit_vector (0 to 31);
	B : in bit_vector (0 to 31);
	CinS : in bit;
	S : out bit_vector (0 to 31);
	CoutS : out bit
);
END Somador32Bits;
architecture comportamento of Somador32Bits is  
	signal TempC: bit_vector (0 to 30);
component manchester
PORT (
	A, B, Cin: in bit;
	S, Cout : out bit
);
end component;
BEGIN 
	m1: manchester
		port map(A => A(0), B => B(0), S => S(0), Cin => CinS, Cout => TempC(0));
	m2: manchester
		port map(A => A(1), B => B(1), S => S(1), Cin => TempC(0), Cout => TempC(1));
	m3: manchester
		port map(A => A(2), B => B(2), S => S(2), Cin => TempC(1), Cout => TempC(2));
	m4: manchester
		port map(A => A(3), B => B(3), S => S(3), Cin => TempC(2), Cout => TempC(3));
	m5: manchester
		port map(A => A(4), B => B(4), S => S(4), Cin => TempC(3), Cout => TempC(4));
	m6: manchester
		port map(A => A(5), B => B(5), S => S(5), Cin => TempC(4), Cout => TempC(5));
	m7: manchester
		port map(A => A(6), B => B(6), S => S(6), Cin => TempC(5), Cout => TempC(6));
	m8: manchester
		port map(A => A(7), B => B(7), S => S(7), Cin => TempC(6), Cout => TempC(7));
	m9: manchester
		port map(A => A(8), B => B(8), S => S(8), Cin => TempC(7), Cout => TempC(8));
	m10: manchester
		port map(A => A(9), B => B(9), S => S(9), Cin => TempC(8), Cout => TempC(9));
	m11: manchester
		port map(A => A(10), B => B(10), S => S(10), Cin => TempC(9), Cout => TempC(10));
	m12: manchester
		port map(A => A(11), B => B(11), S => S(11), Cin => TempC(10), Cout => TempC(11));
	m13: manchester
		port map(A => A(12), B => B(12), S => S(12), Cin => TempC(11), Cout => TempC(12));
	m14: manchester
		port map(A => A(13), B => B(13), S => S(13), Cin => TempC(12), Cout => TempC(13));
	m15: manchester
		port map(A => A(14), B => B(14), S => S(14), Cin => TempC(13), Cout => TempC(14));
	m16: manchester
		port map(A => A(15), B => B(15), S => S(15), Cin => TempC(14), Cout => TempC(15));
	m17: manchester
		port map(A => A(16), B => B(16), S => S(16), Cin => TempC(15), Cout => TempC(16));
	m18: manchester
		port map(A => A(17), B => B(17), S => S(17), Cin => TempC(16), Cout => TempC(17));
	m19: manchester
		port map(A => A(18), B => B(18), S => S(18), Cin => TempC(17), Cout => TempC(18));
	m20: manchester
		port map(A => A(19), B => B(19), S => S(19), Cin => TempC(18), Cout => TempC(19));
	m21: manchester
		port map(A => A(20), B => B(20), S => S(20), Cin => TempC(19), Cout => TempC(20));
	m22: manchester
		port map(A => A(21), B => B(21), S => S(21), Cin => TempC(20), Cout => TempC(21));
	m23: manchester
		port map(A => A(22), B => B(22), S => S(22), Cin => TempC(21), Cout => TempC(22));
	m24: manchester
		port map(A => A(23), B => B(23), S => S(23), Cin => TempC(22), Cout => TempC(23));
	m25: manchester
		port map(A => A(24), B => B(24), S => S(24), Cin => TempC(23), Cout => TempC(24));
	m26: manchester
		port map(A => A(25), B => B(25), S => S(25), Cin => TempC(24), Cout => TempC(25));
	m27: manchester
		port map(A => A(26), B => B(26), S => S(26), Cin => TempC(25), Cout => TempC(26));
	m28: manchester
		port map(A => A(27), B => B(27), S => S(27), Cin => TempC(26), Cout => TempC(27));
	m29: manchester
		port map(A => A(28), B => B(28), S => S(28), Cin => TempC(27), Cout => TempC(28));
	m30: manchester
		port map(A => A(29), B => B(29), S => S(29), Cin => TempC(28), Cout => TempC(29));
	m31: manchester
		port map(A => A(30), B => B(30), S => S(30), Cin => TempC(29), Cout => TempC(30));
	m32: manchester
		port map(A => A(31), B => B(31), S => S(31), Cin => TempC(30), Cout => CoutS);
		
end comportamento;